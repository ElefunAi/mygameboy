// ほぼ未メンテ, 変更行にはGコメあり

`include "define.vh"
module DECODER (
    input wire [7:0] inst, //G
    output wire [31:0] imm,
    output wire [4:0] rs1_addr, rs2_addr, rd_addr,
    output wire [4:0] exe_fun,
    output wire mem_wen, rf_wen,
    output wire [1:0] rs1, wb_sel,
    output wire [2:0] rs2
);
    // 宣言
    // G 内部信号 
    wire [7:0] opcode;
    // wire [4:0] rd;

    // assign
    assign opcode = inst[7:0];
    // デコーダが渡すもの
    // G 16bit長命令ではaluにstall渡してalu側にnop実行してもらう

    // exe_fun(演算内容),rs1(第1オペランド),rs2(第2オペランド),mem_wen(メモリenable),
    // rf_wen(ライトバックenable),wb_sel(ライトバックデータセレクタ)
    // wb_selで例えばWB_ALUは、ALUの出力をレジスタへ書き戻すことを表す
    // つまり、reg_fileにとってはWB_ALU & rf_wen(Write ENable)がenable信号
    // reg_fileに対して=>32bit rs1_addr, rs2_addr, rd_addr, imm(即値)
    assign rs1_addr = inst[19:15];
    assign rs2_addr = inst[24:20];
    assign rd_addr = inst[11:7];
    // 即値の扱い方 risc-v ISA manual参照(P.24)
    assign imm = (opcode == `LUI || opcode == `AUIPC) ? {inst[31:12], 12'd0} : // U-format
                 (opcode == `JAL) ? {{11{inst[31]}},inst[31],inst[19:12],inst[20],inst[30:21],1'd0} : // J-format
                 (opcode == `JALR || opcode == `LW || opcode == `OPIMI) ? {{20{inst[31]}},inst[31],inst[30:25],inst[24:21],inst[20]} : // I-format
                 (opcode == `BRANCH) ? {{19{inst[31]}},inst[31],inst[7],inst[30:25],inst[11:8],1'd0} : //B-format
                 (opcode == `STORE) ? {{20{inst[31]}},inst[31],inst[30:25],inst[11:8],inst[7]} : 32'd0;// ? S-format : R-format(即値なし)

    // G マシンサイクルが命令ごとに異なるので、解釈のためのFFを自分で持つ

    function [7:0] decode;
        input [7:0] opcode;
        if (opcode == `CB) begin
            cb_decode(opcode);
        end

        case (opcode)
            8'h0 :  ports = {`ALU_X, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // NOP    
            8'h10 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // STOP   
            8'h20 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // JR_NZ  
            8'h30 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // JR_NC  
            8'h01 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_BC
            8'h11 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_DE
            8'h21 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_HL
            8'h31 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_SP
            8'h02 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD_BC  
            8'h12 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD_DE  
            8'h22 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD_HLI 
            8'h32 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD_HLD 
            8'h03 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // INC16_BC  
            8'h13 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // INC16_DE
            8'h23 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // INC16_HL  
            8'h33 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // INC16_SP  
            8'h04 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_BC
            8'h14 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_DE
            8'h24 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_HL
            8'h34 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // LD16_SP
            8'h05 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h15 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h25 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h35 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h06 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h16 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h26 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h36 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h07 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h17 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h27 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h37 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h08 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h18 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h28 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h38 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h09 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h19 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h29 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h39 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h40 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h50 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h60 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h70 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h41 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h51 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h61 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h71 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h42 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h52 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h62 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h72 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h43 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h53 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h63 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h73 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h44 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h54 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h64 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h74 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h45 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h55 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h65 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h75 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h46 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h56 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h66 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h76 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h47 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h57 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h67 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h77 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h48 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h58 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h68 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h78 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h49 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h59 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h69 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h79 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h80 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h90 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h81 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h91 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h82 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h92 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h83 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h93 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h84 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h94 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h85 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h95 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h86 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h96 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h87 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h97 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h88 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h98 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h89 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h99 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hED : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            default: begin //NOP=>_Xで統一 
                ports = {`ALU_X, `RS1_X, `RS2_X, `MEN_X, `REN_X, `WB_X};
            end
        endcase       
    endfunction

    // prefix cbの呼び出し
    function cb_decode;
        case (opcode)
            8'h0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU};  // 
            8'h10 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h20 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h30 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h01 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h11 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h21 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h31 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h02 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h12 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h22 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h32 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h03 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h13 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h23 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h33 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h04 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h14 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h24 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h34 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h05 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h15 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h25 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h35 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h06 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h16 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h26 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h36 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h07 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h17 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h27 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h37 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h08 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h18 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h28 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h38 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h09 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h19 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h29 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h39 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h0F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h1F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h2F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h3F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h40 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h50 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h60 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h70 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h41 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h51 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h61 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h71 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h42 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h52 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h62 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h72 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h43 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h53 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h63 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h73 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h44 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h54 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h64 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h74 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h45 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h55 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h65 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h75 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h46 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h56 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h66 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h76 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h47 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h57 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h67 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h77 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h48 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h58 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h68 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h78 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h49 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h59 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h69 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h79 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h4F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h5F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h6F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h7F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h80 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h90 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h81 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h91 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h82 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h92 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h83 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h93 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h84 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h94 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h85 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h95 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h86 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h96 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h87 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h97 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h88 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h98 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h89 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h99 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hA9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hB9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9A : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9B : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9C : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9D : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9E : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h8F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'h9F : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hAF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hBF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF0 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF1 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF2 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF3 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF4 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF5 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF6 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF7 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF8 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hC9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hD9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hE9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hF9 : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFA : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFB : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFC : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hED : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFD : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFE : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hCF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hDF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hEF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            8'hFF : ports = {`ALU_ADD, `RS1_X, `RS2_IMI, `MEN_X, `REN_S, `WB_ALU}; // 
            default: 
        endcase
    endfunction
    
    wire [13:0] probe;
    assign probe = ports(opcode, funct3, funct7);
    assign {exe_fun, rs1, rs2, mem_wen, rf_wen, wb_sel} = ports(opcode, funct3, funct7);
endmodule